module moduleName (
    
);
    
endmodule