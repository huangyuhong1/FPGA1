module key_beep (
    input clk,rst_n
);
    
endmodule